//这是一个非门
module top{
    input in;
    output out;
}

assign out = ~in;

endmodule