module notLatch(
    input in,
    output out);
    
    assign out = ~in;

endmodule
